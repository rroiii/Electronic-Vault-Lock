library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity password_decrypter is
    port (
        encrypted_password : in STD_LOGIC_VECTOR (11 downto 0);
        encrypted_password : out STD_LOGIC_VECTOR (11 downto 0)
    );
end entity password_decrypter;

architecture rtl of password_decrypter is
    
begin
    
    
    
end architecture rtl;